`ifndef __HW_INFO_H__
`define __HW_INFO_H__


`define PLATFORM_ADDR 32
`define NUM_CORE_USER 1
`define NUM_CORE_TEAM 1
`define NUM_LOCK_USER 0
`define NUM_LOCK_SYSTEM 0
`define NUM_BARRIER_USER 0
`define NUM_BARRIER_SYSTEM 0
`define NUM_AUTO_ID 0
`define NUM_GLOBAL_TAG 0
`define SRAM_SIZE (32'h 20000)
`define SRAM_CELL_SIZE (32'h 20000)
`define SRAM_CELL_WIDTH 32
`define SRAM_PORT_WIDTH 32
`define INCLUDE_IROM
`define TICK_HZ 1000000
`define SYSTEM_CLK_HZ 50000000
`define CORE_CLK_HZ 50000000
`define UART_CLK_HZ 50000000
`define SPI_CLK_HZ 50000000
`define I2C_CLK_HZ 50000000
`define OLED_CLK_HZ 50000000
`define PACT_CLK_HZ 0
`define NUM_UART_READYMADE 0
`define NUM_SPI_READYMADE 0
`define NUM_I2C_READYMADE 0
`define NUM_UART_USER 0
`define NUM_SPI_USER 0
`define NUM_I2C_USER 0
`define NUM_LED_CHECKER 0
`define NUM_AIOIF 0
`define NUM_SWITCH_SLIDE_READYMADE 0
//`define INCLUDE_SLOW_DRAM
//`define INCLUDE_FAST_DRAM
//`define INCLUDE_SDRAM
//`define INCLUDE_EXT_MRAM
//`define INCLUDE_DDR
`define INCLUDE_SMALL_RAM
//`define INCLUDE_LARGE_RAM
//`define INCLUDE_BOOT_MODE
//`define INCLUDE_CACHE
//`define INCLUDE_TIMER
//`define INCLUDE_PLIC
//`define INCLUDE_CORE_JTAG
//`define INCLUDE_OLED
//`define INCLUDE_OLED_BW
//`define INCLUDE_OLED_RGB
//`define INCLUDE_SPI_FLASH
`define INCLUDE_UART_PRINTF
//`define INCLUDE_OLEDBW_PRINTF
//`define INCLUDE_FUSE_BOX
//`define INCLUDE_ADC
//`define INCLUDE_USER_INTERRUPTS
//`define INCLUDE_ARDUCAM
//`define INCLUDE_BLUETOOTH
//`define INCLUDE_WIFI
//`define INCLUDE_JPEG_ENCODER
//`define INCLUDE_JPEGLS_ENCODER
//`define INCLUDE_HBC1_TX
//`define INCLUDE_HBC1_RX
//`define INCLUDE_HBC1
`define INCLUDE_CORE_PERI_GROUP
//`define INCLUDE_NOC_DEBUG
//`define INCLUDE_PACT
//`define INCLUDE_STARC
//`define INCLUDE_DCA
//`define INCLUDE_I2S
//`define INCLUDE_DMA
//`define INCLUDE_FLORIAN
//`define INCLUDE_FLORIAN_SP
//`define INCLUDE_FLORIAN_DP
//`define INCLUDE_TRAFFIC_GENERATOR
//`define INCLUDE_VTA
//`define INCLUDE_LCD_SHIELD
//`define INCLUDE_GPIO_PINMUX
//`define INCLUDE_USER_DDR4
//`define INCLUDE_USER_DDR3
//`define INCLUDE_C2C
//`define INCLUDE_EXTINPUT_BACKEND
//`define INCLUDE_EDGE_VIDEO_SYSTEM
//`define INCLUDE_VDMA
//`define INCLUDE_VIM
//`define INCLUDE_VOM
//`define INCLUDE_HDMI
//`define INCLUDE_CIS
//`define INCLUDE_SPI_LCD
//`define INCLUDE_TFT_LCD
//`define INCLUDE_TCACHING
//`define INCLUDE_HW_BARRIER
//`define I2S_SAMPLING_RATE
//`define I2S_IP_CLK_HZ
//`define I2S_MCLK_HZ
`define NOC_FLIT_DIVISOR 1
`define NUM_TRAFFIC_GENERATOR 0
`define NUM_VTA 0
`define NUM_C2C_MASTER 0
`define NUM_C2C_SLAVE 0
`define FIXED_CACHEABLE_START (32'h 00000000)
`define FIXED_CACHEABLE_LAST (32'h bfffffff)
`define PLATFORM_NAME "test_prj_mj2"
`define INCLUDE_RVC_ORCA
`define NUM_CORE 1
`define NUM_REAL_CORE 1
//`define INCLUDE_MULTICORE
`define NUM_BARRIER 0
`define NUM_LOCK 0
`define SPI_INDEX_FOR_READYMADE 0
`define SPI_INDEX_FOR_USER 0
`define SPI_INDEX_FOR_SYSTEM 0
`define NUM_SPI_SYSTEM 0
`define UART_INDEX_FOR_READYMADE 0
`define UART_INDEX_FOR_USER 0
`define UART_INDEX_FOR_SYSTEM 0
`define UART_INDEX_FOR_UART_PRINTF 0
`define NUM_UART_SYSTEM 1
`define I2C_INDEX_FOR_READYMADE 0
`define I2C_INDEX_FOR_USER 0
`define I2C_INDEX_FOR_SYSTEM 0
`define NUM_I2C_SYSTEM 0
`define NUM_GPIO 0
`define NUM_UART 1
`define NUM_SPI 0
`define NUM_I2C 0
`define INCLUDE_CORE_USER
`define INCLUDE_CORE_TEAM
//`define INCLUDE_LOCK_USER
//`define INCLUDE_LOCK_SYSTEM
//`define INCLUDE_BARRIER_USER
//`define INCLUDE_BARRIER_SYSTEM
//`define INCLUDE_AUTO_ID
//`define INCLUDE_GLOBAL_TAG
//`define INCLUDE_UART_READYMADE
//`define INCLUDE_SPI_READYMADE
//`define INCLUDE_I2C_READYMADE
//`define INCLUDE_UART_USER
//`define INCLUDE_SPI_USER
//`define INCLUDE_I2C_USER
//`define INCLUDE_LED_CHECKER
//`define INCLUDE_AIOIF
//`define INCLUDE_SWITCH_SLIDE_READYMADE
//`define INCLUDE_C2C_MASTER
//`define INCLUDE_C2C_SLAVE
`define INCLUDE_CORE
`define INCLUDE_REAL_CORE
//`define INCLUDE_BARRIER
//`define INCLUDE_LOCK
//`define INCLUDE_SPI_SYSTEM
`define INCLUDE_UART_SYSTEM
//`define INCLUDE_I2C_SYSTEM
//`define INCLUDE_GPIO
`define INCLUDE_UART
//`define INCLUDE_SPI
//`define INCLUDE_I2C
`define NUM_PREDEFINED_CLOCK 0
`define INCLUDE_SRAM
//`define INCLUDE_DRAM

`endif
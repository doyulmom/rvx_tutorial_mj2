wire [BW_USERNAME-1:0] username_string = `FORMAT_STRING("None");
wire [BW_GIT_NAME-1:0] home_git_name_string = `FORMAT_STRING("rvx_tutorial_mj2");
wire [BW_GIT_VERSION-1:0] home_git_version_string = `FORMAT_STRING("cfc87d6");
wire [BW_GIT_VERSION-1:0] devkit_git_version_string = `FORMAT_STRING("fc2cb49");
wire [BW_DATE-1:0] design_date_string = `FORMAT_STRING("2025-08-08 11:21");